module test ();

    $display("hello,world");
    
endmodule